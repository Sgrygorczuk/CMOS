*** SPICE deck for cell nmos_iv{sch} from library tutorial_2
*** Created on Mon Feb 18, 2019 13:10:11
*** Last revised on Mon Feb 18, 2019 15:06:05
*** Written on Mon Feb 18, 2019 15:06:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd

*** TOP LEVEL CELL: nmos_iv{sch}
Mnmos-4@0 d g s gnd NMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'nmos_iv{sch}'
vs s 0 DC 0
vw w 0 DC 0 
vg g 0 DC 0
vd d 0 dC 0
.dc vd 0 5 1m vg 0 5 1  
.include D:\Programs\Electric\C5_models.txt
.END
