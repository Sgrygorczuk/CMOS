* First line is ignored

*** SUBCIRCUIT TEEST FROM CELL TEEST{lay}
.SUBCKT TEEST gnd Out_1 Out_2 Out_3 vdd X Y
Mnmos@0 Out_2 X gnd gnd N L=0.7U W=1.75U
Mnmos@1 Out_1 Y gnd gnd N L=0.7U W=1.75U
Mnmos@2 net@80 Out_1 gnd gnd N L=0.7U W=1.75U
Mnmos@3 gnd Y net@101 gnd N L=0.7U W=1.75U
Mnmos@4 net@101 Out_2 Out_3 gnd N L=0.7U W=1.75U
Mnmos@5 Out_3 X net@80 gnd N L=0.7U W=1.75U
Mpmos@0 Out_2 X vdd vdd P L=0.7U W=1.75U
Mpmos@1 Out_1 Y vdd vdd P L=0.7U W=1.75U
Mpmos@2 net@200 Out_1 vdd vdd P L=0.7U W=1.75U
Mpmos@3 Out_3 Y net@200 vdd P L=0.7U W=1.75U
Mpmos@4 vdd X net@200 vdd P L=0.7U W=1.75U
Mpmos@6 net@200 Out_2 Out_3 vdd P L=0.7U W=1.75U
.ENDS TEEST
