*** SPICE deck for cell 32_Adder{lay} from library Project_3
*** Created on Sat May 11, 2019 23:57:42
*** Last revised on Sun May 12, 2019 18:43:08
*** Written on Sun May 12, 2019 18:43:30 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project_3__Full_Adder FROM CELL Full_Adder{lay}
.SUBCKT Project_3__Full_Adder A B C C0 G gnd P S vdd
Mnmos@21 net@369 net@353 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=3.828P PS=24.35U PD=7.875U
Mnmos@22 gnd B net@388 gnd N L=0.7U W=1.75U AS=1.531P AD=16.713P PS=3.5U PD=24.35U
Mnmos@23 net@388 C0 net@390 gnd N L=0.7U W=1.75U AS=2.527P AD=1.531P PS=4.637U PD=3.5U
Mnmos@24 net@390 net@358 net@369 gnd N L=0.7U W=1.75U AS=3.828P AD=2.527P PS=7.875U PD=4.637U
Mnmos@25 net@358 C0 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.288P PS=24.35U PD=8.4U
Mnmos@26 net@353 B gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.441P PS=24.35U PD=8.575U
Mnmos@27 net@461 net@445 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=3.828P PS=24.35U PD=7.875U
Mnmos@28 gnd A net@480 gnd N L=0.7U W=1.75U AS=1.531P AD=16.713P PS=3.5U PD=24.35U
Mnmos@29 net@480 net@390 P gnd N L=0.7U W=1.75U AS=2.527P AD=1.531P PS=4.637U PD=3.5U
Mnmos@30 P net@450 net@461 gnd N L=0.7U W=1.75U AS=3.828P AD=2.527P PS=7.875U PD=4.637U
Mnmos@31 net@450 net@390 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.594P PS=24.35U PD=8.75U
Mnmos@32 net@445 A gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.441P PS=24.35U PD=8.575U
Mnmos@33 net@553 net@537 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=3.828P PS=24.35U PD=7.875U
Mnmos@34 gnd C net@572 gnd N L=0.7U W=1.75U AS=1.531P AD=16.713P PS=3.5U PD=24.35U
Mnmos@35 net@572 P S gnd N L=0.7U W=1.75U AS=2.527P AD=1.531P PS=4.637U PD=3.5U
Mnmos@36 S net@542 net@553 gnd N L=0.7U W=1.75U AS=3.828P AD=2.527P PS=7.875U PD=4.637U
Mnmos@37 net@542 P gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.288P PS=24.35U PD=8.4U
Mnmos@38 net@537 C gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.441P PS=24.35U PD=8.575U
Mnmos@39 gnd net@390 net@654 gnd N L=0.7U W=1.75U AS=3.369P AD=16.713P PS=5.6U PD=24.35U
Mnmos@40 net@654 A net@645 gnd N L=0.7U W=1.75U AS=3.879P AD=3.369P PS=6.767U PD=5.6U
Mnmos@41 G net@645 gnd gnd N L=0.7U W=1.75U AS=16.713P AD=4.288P PS=24.35U PD=8.4U
Mpmos@21 net@352 net@353 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=2.909P PS=25.247U PD=5.075U
Mpmos@22 vdd net@358 net@352 vdd P L=0.7U W=1.75U AS=2.909P AD=16.823P PS=5.075U PD=25.247U
Mpmos@23 net@390 B net@352 vdd P L=0.7U W=1.75U AS=2.909P AD=2.527P PS=5.075U PD=4.637U
Mpmos@24 net@352 C0 net@390 vdd P L=0.7U W=1.75U AS=2.527P AD=2.909P PS=4.637U PD=5.075U
Mpmos@25 net@358 C0 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.288P PS=25.247U PD=8.4U
Mpmos@26 net@353 B vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.441P PS=25.247U PD=8.575U
Mpmos@27 net@444 net@445 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=2.909P PS=25.247U PD=5.075U
Mpmos@28 vdd net@450 net@444 vdd P L=0.7U W=1.75U AS=2.909P AD=16.823P PS=5.075U PD=25.247U
Mpmos@29 P A net@444 vdd P L=0.7U W=1.75U AS=2.909P AD=2.527P PS=5.075U PD=4.637U
Mpmos@30 net@444 net@390 P vdd P L=0.7U W=1.75U AS=2.527P AD=2.909P PS=4.637U PD=5.075U
Mpmos@31 net@450 net@390 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.594P PS=25.247U PD=8.75U
Mpmos@32 net@445 A vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.441P PS=25.247U PD=8.575U
Mpmos@33 net@536 net@537 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=2.909P PS=25.247U PD=5.075U
Mpmos@34 vdd net@542 net@536 vdd P L=0.7U W=1.75U AS=2.909P AD=16.823P PS=5.075U PD=25.247U
Mpmos@35 S C net@536 vdd P L=0.7U W=1.75U AS=2.909P AD=2.527P PS=5.075U PD=4.637U
Mpmos@36 net@536 P S vdd P L=0.7U W=1.75U AS=2.527P AD=2.909P PS=4.637U PD=5.075U
Mpmos@37 net@542 P vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.288P PS=25.247U PD=8.4U
Mpmos@38 net@537 C vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.441P PS=25.247U PD=8.575U
Mpmos@39 vdd net@390 net@645 vdd P L=0.7U W=1.75U AS=3.879P AD=16.823P PS=6.767U PD=25.247U
Mpmos@40 net@645 A vdd vdd P L=0.7U W=1.75U AS=16.823P AD=3.879P PS=25.247U PD=6.767U
Mpmos@41 G net@645 vdd vdd P L=0.7U W=1.75U AS=16.823P AD=4.288P PS=25.247U PD=8.4U
.ENDS Project_3__Full_Adder

*** TOP LEVEL CELL: 32_Adder{lay}
XFull_Add@0 A0 B0 C0 C0 G0 gnd P0 S0 vdd Project_3__Full_Adder
XFull_Add@1 A1 B1 C1 C0 G1 gnd P1 S1 vdd Project_3__Full_Adder
XFull_Add@2 A2 B2 C2 C0 G2 gnd P2 S2 vdd Project_3__Full_Adder
XFull_Add@3 A3 B3 C3 C0 G3 gnd P3 S3 vdd Project_3__Full_Adder
XFull_Add@4 A4 B4 C4 C0 G4 gnd P4 S4 vdd Project_3__Full_Adder
XFull_Add@5 A5 B5 C5 C0 G5 gnd P5 S5 vdd Project_3__Full_Adder
XFull_Add@6 A6 B6 C6 C0 G6 gnd P6 S6 vdd Project_3__Full_Adder
XFull_Add@7 A7 B7 C7 C0 G7 gnd P7 S7 vdd Project_3__Full_Adder
XFull_Add@8 A8 B8 C8 C0 G8 gnd P8 S8 vdd Project_3__Full_Adder
XFull_Add@9 A9 B9 C9 C0 G9 gnd P9 S9 vdd Project_3__Full_Adder
XFull_Add@10 A10 B10 C10 C0 G10 gnd P10 S10 vdd Project_3__Full_Adder
XFull_Add@11 A11 B11 C11 C0 G11 gnd P11 S11 vdd Project_3__Full_Adder
XFull_Add@12 A12 B12 C12 C0 G12 gnd P12 S12 vdd Project_3__Full_Adder
XFull_Add@13 A13 B13 C13 C0 G13 gnd P13 S13 vdd Project_3__Full_Adder
XFull_Add@14 A14 B14 C14 C0 G14 gnd P14 S14 vdd Project_3__Full_Adder
XFull_Add@15 A15 B15 C15 C0 G15 gnd P15 S15 vdd Project_3__Full_Adder
XFull_Add@16 A16 B16 C16 C0 G16 gnd P16 S16 vdd Project_3__Full_Adder
XFull_Add@17 A17 B17 C17 C0 G17 gnd P17 S17 vdd Project_3__Full_Adder
XFull_Add@18 A18 B18 C18 C0 G18 gnd P18 S18 vdd Project_3__Full_Adder
XFull_Add@19 A19 B19 C19 C0 G19 gnd P19 S19 vdd Project_3__Full_Adder
XFull_Add@20 A20 B20 C20 C0 G20 gnd P20 S20 vdd Project_3__Full_Adder
XFull_Add@21 A21 B21 C21 C0 G21 gnd P21 S21 vdd Project_3__Full_Adder
XFull_Add@22 A22 B22 C22 C0 G22 gnd P22 S22 vdd Project_3__Full_Adder
XFull_Add@23 A23 B23 C23 C0 G23 gnd P23 S23 vdd Project_3__Full_Adder
XFull_Add@24 A24 B24 C24 C0 G24 gnd P24 S24 vdd Project_3__Full_Adder
XFull_Add@25 A25 B25 C25 C0 G25 gnd P25 S25 vdd Project_3__Full_Adder
XFull_Add@26 A26 B26 C26 C0 G26 gnd P26 S26 vdd Project_3__Full_Adder
XFull_Add@27 A27 B27 C27 C0 G27 gnd P27 S27 vdd Project_3__Full_Adder
XFull_Add@28 A28 B28 C28 C0 G28 gnd P28 S28 vdd Project_3__Full_Adder
XFull_Add@29 A29 B29 C29 C0 G29 gnd P29 S29 vdd Project_3__Full_Adder
XFull_Add@30 A30 B30 C30 C0 G30 gnd P30 S30 vdd Project_3__Full_Adder
XFull_Add@31 A31 B31 C31 C0 G31 gnd P31 S31 vdd Project_3__Full_Adder

* Spice Code nodes in cell cell '32_Adder{lay}'
VDD VDD 0 DC 3.3 
VGND GND 0 DC 0
VIN2 A0 0 PULSE(3.3 0 0 1n 1n 20n 40n)
VIN3 A1 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN4 A2 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN5 A3 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN6 A4 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN7 A5 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN8 A6 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN9 A7 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN10 A8 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN11 A9 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN12 A10 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN13 A11 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN14 A12 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN15 A13 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN16 A14 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN17 A15 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN18 A16 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN19 A17 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN20 A18 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN21 A19 0 PULSE(3.3 0 0 1n 1n 160n 320n
VIN22 A20 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN23 A21 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN24 A22 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN25 A23 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN26 A24 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN27 A25 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN28 A26 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN29 A27 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN30 A28 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN31 A29 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN32 A30 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN33 A31 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN97 B0 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN34 B1 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN35 B2 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN36 B3 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN37 B4 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN38 B5 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN39 B6 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN40 B7 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN41 B8 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN42 B9 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN43 B10 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN44 B11 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN45 B12 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN46 B13 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN47 B14 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN48 B15 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN49 B16 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN50 B17 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN51 B18 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN52 B19 0 PULSE(3.3 0 0 1n 1n 160n 320n
VIN53 B20 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN54 B21 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN55 B22 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN56 B23 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN57 B24 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN58 B25 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN59 B26 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN60 B27 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN61 B28 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN62 B29 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN63 B30 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN64 B31 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN65 C0 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN66 C1 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN67 C2 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN68 C3 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN69 C4 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN70 C5 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN71 C6 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN72 C7 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN73 C8 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN74 C9 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN75 C10 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN76 C11 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN77 C12 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN78 C13 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN79 C14 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN80 C15 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN81 C16 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN82 C17 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN83 C18 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN84 C19 0 PULSE(3.3 0 0 1n 1n 160n 320n
VIN85 C20 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN86 C21 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN87 C22 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN88 C23 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN89 C24 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN90 C25 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN91 C26 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN92 C27 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN93 C28 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN94 C29 0  PULSE(3.3 0 0 1n 1n 160n 320n)
VIN95 C30 0 PULSE(3.3 0 0 1n 1n 160n 320n)
VIN96 C31 0 PULSE(3.3 0 0 1n 1n 160n 320n)
.TRAN 0 59n
.include C:\electric\MOS_model.txt
.END
