*** SPICE deck for cell XOR_PART_1{lay} from library Project-2
*** Created on Sat Apr 06, 2019 19:57:40
*** Last revised on Sat Apr 06, 2019 20:00:36
*** Written on Sun Apr 07, 2019 13:47:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: XOR_PART_1{lay}
Mnmos@0 net@27 D gnd gnd N L=0.7U W=1.75U AS=14.547P AD=3.981P PS=20.125U PD=8.05U
Mnmos@1 gnd B net@41 gnd N L=0.7U W=1.75U AS=1.531P AD=14.547P PS=3.5U PD=20.125U
Mnmos@2 net@41 A F gnd N L=0.7U W=1.75U AS=2.45P AD=1.531P PS=4.55U PD=3.5U
Mnmos@3 F C net@27 gnd N L=0.7U W=1.75U AS=3.981P AD=2.45P PS=8.05U PD=4.55U
Mpmos@0 net@0 D vdd vdd P L=0.7U W=1.75U AS=16.231P AD=2.909P PS=25.55U PD=5.075U
Mpmos@1 vdd C net@0 vdd P L=0.7U W=1.75U AS=2.909P AD=16.231P PS=5.075U PD=25.55U
Mpmos@2 F B net@0 vdd P L=0.7U W=1.75U AS=2.909P AD=2.45P PS=5.075U PD=4.55U
Mpmos@3 net@0 A F vdd P L=0.7U W=1.75U AS=2.45P AD=2.909P PS=4.55U PD=5.075U

* Spice Code nodes in cell cell 'XOR_PART_1{lay}'
VDD VDD 0 DC 3.3 
VGND GND 0 DC 0
VIN A 0 PULSE(3.3 0 0 100p 100p 10n 20n)
VIN2 B 0 PULSE(3.3 0 0 100p 100p 20n 40n)
VIN3 C 0 PULSE(0 3.3 0 100p 100p 10n 20n)
VIN4 D 0 PULSE(0 3.3 0 100p 100p 20n 40n)
.TRAN 0 40n
.include C:\electric\MOS_model.txt
.END
