*** SPICE deck for cell inv_20_10{sch} from library tutorial_3
*** Created on Mon Feb 18, 2019 16:23:34
*** Last revised on Tue Feb 19, 2019 18:07:20
*** Written on Tue Feb 19, 2019 18:14:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inv_20_10{sch}
Mnmos-4@0 out in gnd gnd N L=0.7U W=1.4U
Mpmos-4@0 out in vdd vdd P L=0.7U W=2.8U

* Spice Code nodes in cell cell 'inv_20_10{sch}'
VDD VDD 0 DC 3.3 
VGND GND 0 DC 0
VIN In 0 PULSE(3.3 0 0 100p 100p 10n 20n)
.TRAN 0 50n
.include D:\Programs\Electric\MOS_model.txt
.END
