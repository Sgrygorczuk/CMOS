*** SPICE deck for cell HW4{lay} from library HW4
*** Created on Mon Apr 29, 2019 09:08:47
*** Last revised on Mon Apr 29, 2019 10:04:09
*** Written on Mon Apr 29, 2019 10:04:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: HW4:HW4{lay}
Mnmos@0 gnd clk F gnd N L=0.7U W=1.75U AS=3.879P AD=53.9P PS=6.767U PD=68.6U
Mnmos@1 F w net@1 gnd N L=0.7U W=1.75U AS=1.838P AD=3.879P PS=3.85U PD=6.767U
Mnmos@2 net@1 x net@4 gnd N L=0.7U W=1.75U AS=1.838P AD=1.838P PS=3.85U PD=3.85U
Mnmos@3 net@4 x net@6 gnd N L=0.7U W=1.75U AS=1.838P AD=1.838P PS=3.85U PD=3.85U
Mnmos@4 F y net@9 gnd N L=0.7U W=1.75U AS=1.838P AD=3.879P PS=3.85U PD=6.767U
Mnmos@5 net@6 z F gnd N L=0.7U W=1.75U AS=3.879P AD=1.838P PS=6.767U PD=3.85U
Mnmos@6 net@9 x F gnd N L=0.7U W=1.75U AS=3.879P AD=1.838P PS=6.767U PD=3.85U
Mpmos@0 vdd clk F vdd P L=0.7U W=1.75U AS=3.879P AD=17.15P PS=6.767U PD=26.6U

* Spice Code nodes in cell cell 'HW4:HW4{lay}'
VDD VDD 0 DC 3.3 
VGND GND 0 DC 0
VIN clk 0 PULSE(3.3 0 0 100p 100p 500p 1000p)
VDD2 x VDD 0 DC 3.3
VIN2 y 0 PULSE(3.3 0 0 100p 100p  2n 4n)
VDD3 w VDD 0 DC 3.3)
VDD4 z VDD 0 DC 3.3
.TRAN 0 12n
.include C:\electric\MOS_model.txt
.END
